module register_controller(


);


endmodule
