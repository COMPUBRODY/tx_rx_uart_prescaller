module register_controller(
			input clock,
			input [7:0] rx_in,
			output [7:0] tx_out,
			output [3:0] Byte_0,
			output [3:0] Byte_1,
			output [3:0] Byte_2,
			output [3:0] Byte_3,
			output [3:0] Byte_4,
			output [3:0] Byte_5
		
);


endmodule
