`timescale 1ns / 10ps

module tb_preescaller();

    reg clock,
    wire enable_flag;




endmodule